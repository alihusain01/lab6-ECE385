
module lab61soc (
	clk_clk,
	reset_reset_n,
	led_wire_export);	

	input		clk_clk;
	input		reset_reset_n;
	output	[7:0]	led_wire_export;
endmodule
